module mode2 (in, out1, out2, out3);
	input in;
	output [3:0] out1, out2, out3;
	
	count AAA (in, out1, out2, out3);
endmodule 